*
R3 2 1 {R}
R5 0 2 {R}
R6 0 3 {R}
V1 1 0 {V}
D1 3 2 D
.model D D
.lib /Users/lancemathias/Library/Application Support/LTspice/lib/cmp/standard.dio
.param V=5
.param R=1
.tran	 1
.backanno
.end
